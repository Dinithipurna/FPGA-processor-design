module core_tb();
