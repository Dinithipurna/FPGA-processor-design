module global_var;

	initial begin
	reg Iin=1;
	reg Iout=0;
	reg Din=1;
	reg Dout=0;
	
	end
endmodule
