module char_7_seg(C,display);
S