package mypkg;
	reg ID;
	reg DD;
	
	initial begin
			ID=1;
			DD=1; 
		end
	
endpackage

