`include "define.v"
 

  module Processor(CLK);//,//rst,en,clk_div);


  wire [1:0] MEMCtrl;

  wire [7:0] DAddress,Ddout,IAddress;

  wire [7:0] Ddin,Idin;
 // wire clk_div;

  input CLK;//,rst,en;
 // output clk_div;
 
 // clkdiv clkdiv1(CLK,rst,en,clk_div);
  TopRegisterWrapper TRW1(MEMCtrl,DAddress,Ddout,Ddin,IAddress,Idin,CLK);
 

  IRAM IRAM1(

	.address(IAddress),

	.clock(CLK),

	.data(),

	.wren(1'b0),

	.q(Idin));

	

	DRAM DRAM1(

	.address(DAddress),

	.clock(CLK),

	.data(Ddout),

	.wren(MEMCtrl[0]),

	.q(Ddin));

  


  endmodule

