module check_cp(Wen, BusOut, Clk, RST, INC, dout);
  input Wen, Clk, RST, INC;
  input[3:0] BusOut;
  output reg[3:0] dout = 4'd0;
  reg[3:0] rbase = 4'd0;
  always @(posedge Clk)
    begin
        if (Wen)
            begin
					if((dout == 4'd0))	
					rbase <= BusOut;           
					dout <= BusOut;
            end
        else if (RST) dout <= rbase;
        else if (INC) dout <= dout+1;
        else            dout <= dout;
      
    end
endmodule